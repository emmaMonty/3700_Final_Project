`timescale 1ns/1ps
module audio (

);
endmodule