`timescale 1ns/1ps
module tx_testbench ();
    
endmodule //tx_testbench