`timescale 1ns/1ps
module audio_testbench();

endmodule//testbench